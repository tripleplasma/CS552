module memory_wb_latch(clk, rst, readData_m, readData_wb, aluOut_m, aluOut_wb, memToReg_m, memToReg_wb, link_m, link_wb);

    input wire clk, rst;

endmodule